module covered_vpi;
initial $covered_sim( "delay1.3.cdd", main );
endmodule
